* Resistor Netlist with Sky130 Model

.include /home/monica/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__res_xhigh_po__base.model.spice
.include /home/monica/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__res_xhigh_po_0p35.model.spice

.param sky130_fd_pr__res_high_po__var_mult=1 crpf_precision=1 crpfsw_precision_1_1=1 mc_mm_switch=0

* Instantiate the resistor from top to ground
X0 top 0 0 sky130_fd_pr__res_xhigh_po_0p35 l=1.01 w=0.35 mult=1

* Voltage source
V1 top 0 DC 1

.control
op
print i(V1)
.endc

.end







