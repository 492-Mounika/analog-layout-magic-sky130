* SPICE3 file created for RC circuit with 2fF capacitor - technology: sky130A

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Voltage Source - 1.8V pulse input
V1 IN 0 PULSE(0 1.8 0 100p 100p 1n 10n)

* Resistor - 10kΩ between IN and OUT
R1 IN OUT 10k

* Capacitor instance - 2fF using MIM capacitor (sky130_fd_pr__cap_mim_m3_1)
* Effective capacitance depends on L and W; 1x1 might give ~1fF. Double it for 2fF.
X0 OUT 0 sky130_fd_pr__cap_mim_m3_1 l=2 w=1

.control
tran 1p 20n
plot v(IN) v(OUT)
.endc

.end


