* SPICE3 file created from potentialdiv2.ext - technology: sky130A

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

V1 VDD 0 DC 1.8

* Resistor R1: 3k (shorter length)
X0 VDD OUT GND sky130_fd_pr__res_xhigh_po_0p35 l=0.69

* Resistor R2: 12k (longer length)
X1 OUT GND GND sky130_fd_pr__res_xhigh_po_0p35 l=2.26

.control
tran 1n 10n
print v(OUT)
.endc

.end



